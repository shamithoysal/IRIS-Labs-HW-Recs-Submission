`timescale 1 ns / 1 ps

module dataproc_tb;
    reg clk;
    always #5 clk = (clk === 1'b0);  // 100 MHz

    reg [5:0] reset_cnt = 0;
    wire resetn = &reset_cnt;

    always @(posedge clk) begin
        reset_cnt <= reset_cnt + !resetn;
    end

    localparam ser_half_period = 10;
    event ser_sample;

    wire ser_rx;
    wire ser_tx;

    wire flash_csb;
    wire flash_clk;
    wire flash_io0;
    wire flash_io1;
    wire flash_io2;
    wire flash_io3;

    // Instantiate the SoC wrapper with 128 KB RAM (MEM_WORDS = 32768)
    rvsoc_wrapper #(
        .MEM_WORDS(32768)
    ) uut (
        .clk      (clk),
        .resetn   (resetn),
        .ser_rx   (ser_rx),
        .ser_tx   (ser_tx),
        .flash_csb(flash_csb),
        .flash_clk(flash_clk),
        .flash_io0(flash_io0),
        .flash_io1(flash_io1),
        .flash_io2(flash_io2),
        .flash_io3(flash_io3)
    );

    // External SPI flash model (holds the firmware)
    spiflash spiflash (
        .csb(flash_csb),
        .clk(flash_clk),
        .io0(flash_io0),
        .io1(flash_io1),
        .io2(flash_io2),
        .io3(flash_io3)
    );

    // Load firmware into the flash memory
    initial begin
        $readmemh("firmware.hex", spiflash.memory);
    end

    // Run simulation for 500 us (adjust as needed)
    initial #10000_000 $finish;

    // -----------------------------------------------------------------
    // UART receiver with number accumulation
    // -----------------------------------------------------------------
    reg [7:0] buffer;
    integer current_number;
    reg in_number;

    initial begin
        current_number = 0;
        in_number = 0;
    end

    always begin
        @(negedge ser_tx);

        repeat (ser_half_period) @(posedge clk);
        -> ser_sample;

        repeat (8) begin
            repeat (ser_half_period) @(posedge clk);
            repeat (ser_half_period) @(posedge clk);
            buffer = {ser_tx, buffer[7:1]};
            -> ser_sample;
        end

        repeat (ser_half_period) @(posedge clk);
        repeat (ser_half_period) @(posedge clk);
        -> ser_sample;

        // Process the received character
        if (buffer >= "0" && buffer <= "9") begin
            current_number = current_number * 10 + (buffer - "0");
            in_number = 1;
        end else if (buffer == " " || buffer == "\n" || buffer == "\r") begin
            if (in_number) begin
                $display("Result: %0d", current_number);
                current_number = 0;
                in_number = 0;
            end
        end else begin
            // For other characters (like letters), print them as is
            if (buffer < 32 || buffer >= 127)
                $display("Serial data: %d", buffer);
            else
                $display("Serial data: '%c'", buffer);
        end
    end

    // Optional heartbeat
    always #100_000 $display("[SIM] Time %t", $time);

endmodule